library ieee;
use ieee.std_logic_1164.all;

package ft_pkg is

   type multi32_t is array (integer range <>) of std_logic_vector(31 downto 0);

end package ft_pkg;
