module (		
	input stall
	);
   
      
   default clocking @(posedge clk); endclocking
   default disable iff reset;
   stall_2_clk_max: asse

  
