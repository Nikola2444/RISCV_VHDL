library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity control_path is
  port (clk: in std_logic;
        reset: in std_logic;
        opcode: in std_logic_vector (6 downto 0)
        --***control signal remain to be added***
        
        --***************************************
        );  
end entity;


architecture Behavioral of control_path is
begin
  
end architecture;

