nikola.kovacevic@ws0.lab317.kel.net.3522:1568200739