nikola@nikola.22213:1596270169